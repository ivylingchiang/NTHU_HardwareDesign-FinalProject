module DisplayStack(
  
);

endmodule