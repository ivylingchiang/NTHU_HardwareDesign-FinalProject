module stack(
  input clk,
  input [4:0]state,
  input decision,
  input stackEn,
  output pop,
  output validpop
);
endmodule